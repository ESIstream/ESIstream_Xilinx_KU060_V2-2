-------------------------------------------------------------------------------
-- This is free and unencumbered software released into the public domain.
--
-- Anyone is free to copy, modify, publish, use, compile, sell, or distribute
-- this software, either in source code form or as a compiled bitstream, for 
-- any purpose, commercial or non-commercial, and by any means.
--
-- In jurisdictions that recognize copyright laws, the author or authors of 
-- this software dedicate any and all copyright interest in the software to 
-- the public domain. We make this dedication for the benefit of the public at
-- large and to the detriment of our heirs and successors. We intend this 
-- dedication to be an overt act of relinquishment in perpetuity of all present
-- and future rights to this software under copyright law.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR 
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, 
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN 
-- ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION
-- WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
--
-- THIS DISCLAIMER MUST BE RETAINED AS PART OF THIS FILE AT ALL TIMES. 
-------------------------------------------------------------------------------
-- Version      Date            Author       Description
-- 1.0          2019            Teledyne-e2v Creation
-- 1.1          2019            REFLEXCES    FPGA target migration, 64-bit data path
-- 1.2          2020            Teledyne-e2v Tx emulator, add lss output flag (lane synchronization sequence) 
-------------------------------------------------------------------------------
-- Description :
-- When a sync event occurs, generates the synchronization sequence for receiver frame alignment
-- and PRBS initialization. 
-- Else, 
-- when SER_WIDTH = 32 : it scrambles 2x14-bit ESIstream data with a pseudo-random binary sequence generated by the LFSR module
-- and concatenate the overhead clock bit to each data 
-- when SER_WIDTH = 64 : it scrambles 4x14-bit ESIstream data with a pseudo-random binary sequence generated by the LFSR module
-- and concatenate the overhead clock bit to each data 
----------------------------------------------------------------------------------------------------

library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.esistream_pkg.all;

entity tx_emu_scrambling is
  generic(
    COMMA : std_logic_vector(31 downto 0) := x"FF0000FF"
    );
  port (
    nrst         : in  std_logic;
    clk          : in  std_logic;
    sync         : in  std_logic;                                  -- Start synchronization sequence
    prbs_en      : in  std_logic;                                  -- Enables scrambling processing
    data_in      : in  slv_14_array_n((SER_WIDTH/16)-1 downto 0);  -- Input data to encode
    data_prbs    : in  slv_14_array_n((SER_WIDTH/16)-1 downto 0);
    data_out     : out slv_16_array_n((SER_WIDTH/16)-1 downto 0) := (others => (others => '0'));
    data_out_vld : out std_logic;
    lss          : out std_logic                                   -- when '1' lane synchronization sequence (FAS + PSS) else normal operation.       
    );
end entity tx_emu_scrambling;

architecture rtl of tx_emu_scrambling is
  --============================================================================================================================
  -- Function and Procedure declarations
  --============================================================================================================================

  --============================================================================================================================
  -- Constant and Type declarations
  --============================================================================================================================
  constant NORMAL_OPERATION : std_logic := '0';
  constant SYNC_SEQUENCE    : std_logic := '1';
  constant CLK_BIT_HIGH     : std_logic := '1';
  constant CLK_BIT_LOW      : std_logic := '0';
  --============================================================================================================================
  -- Component declarations
  --============================================================================================================================

  --============================================================================================================================
  -- Signal declarations
  --============================================================================================================================
  signal state    : std_logic                    := '0';  -- '0': NORMAL_OPERATION; '1':SYNC_SEQUENCE
  signal sync_buf : std_logic_vector(1 downto 0) := "00";
  signal cnt_sync : unsigned(4 downto 0)         := (others => '0');
begin
  lss <= state;                                           -- when '1' lane synchronization sequence (FAS + PSS) else normal operation.
  --============================================================================================================================
  -- Sync rising_edge detector
  --============================================================================================================================
  process(clk, nrst)
  begin
    if nrst = '0' then
      sync_buf <= (others => '0');
    elsif rising_edge(clk) then
      sync_buf(0) <= sync;
      sync_buf(1) <= sync_buf(0);
    end if;
  end process;

  --============================================================================================================================
  -- Main FSM
  --============================================================================================================================
  process(clk)
  begin
    if rising_edge(clk) then
      if state = NORMAL_OPERATION then
        cnt_sync                      <= (others => '0');
        data_out_vld                  <= '1';
        if sync_buf = "10" then state <= SYNC_SEQUENCE; data_out_vld <= '0'; end if;
      else  -- SYNC_SEQUENCE 
        cnt_sync                                                  <= cnt_sync + 1;
        if SER_WIDTH = 32 and cnt_sync = 31 then state            <= NORMAL_OPERATION; end if;
        if SER_WIDTH = 32 and cnt_sync(4) = '1' then data_out_vld <= '1'; end if;
        if SER_WIDTH = 64 and cnt_sync = 15 then state            <= NORMAL_OPERATION; end if;
        if SER_WIDTH = 64 and cnt_sync(3) = '1' then data_out_vld <= '1'; end if;
      end if;
    end if;
  end process;

  --============================================================================================================================
  -- Generate the output data according to the FSM and the serialization factor
  --============================================================================================================================
  gen_data_per_ser : for index in 0 to (SER_WIDTH/16)-1 generate
    process(clk)
    begin
      if rising_edge(clk) then
        case (index mod 2) is
          when 0 =>  -- data 0, data 2 (if SER_WIDTH = 32 or 64)
            if state = NORMAL_OPERATION then
              if prbs_en = '1' then data_out(index) <= '0' & CLK_BIT_HIGH & (data_in(index) xor data_prbs(index));
              else data_out(index)                  <= '0' & CLK_BIT_HIGH & data_in(index); end if;
            else     -- SYNC_SEQUENCE
              if SER_WIDTH = 32 and cnt_sync(4) = '0' then data_out(index)                          <= COMMA(15 downto 0);
              elsif SER_WIDTH = 64 and cnt_sync(4) = '0' and cnt_sync(3) = '0' then data_out(index) <= COMMA(15 downto 0);
              else data_out(index)                                                                  <= '0' & CLK_BIT_HIGH & data_prbs(index); end if;
            end if;

          when others =>  -- data 1 (if SER_WIDTH = 32 or 64), data 3 (if SER_WIDTH = 32 or 64)  
            if state = NORMAL_OPERATION then
              if prbs_en = '1' then data_out(index) <= '0' & CLK_BIT_LOW & (data_in(index) xor data_prbs(index));
              else data_out(index)                  <= '0' & CLK_BIT_LOW & data_in(index); end if;
            else          -- SYNC_SEQUENCE   
              if SER_WIDTH = 32 and cnt_sync(4) = '0' then data_out(index)                          <= COMMA(31 downto 16);
              elsif SER_WIDTH = 64 and cnt_sync(4) = '0' and cnt_sync(3) = '0' then data_out(index) <= COMMA(31 downto 16);
              else data_out(index)                                                                  <= '0' & CLK_BIT_LOW & data_prbs(index); end if;
            end if;
        end case;
      end if;
    end process;
  end generate gen_data_per_ser;
end architecture rtl;
