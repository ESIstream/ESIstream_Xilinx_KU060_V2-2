-------------------------------------------------------------------------------
-- This is free and unencumbered software released into the public domain.
--
-- Anyone is free to copy, modify, publish, use, compile, sell, or distribute
-- this software, either in source code form or as a compiled bitstream, for 
-- any purpose, commercial or non-commercial, and by any means.
--
-- In jurisdictions that recognize copyright laws, the author or authors of 
-- this software dedicate any and all copyright interest in the software to 
-- the public domain. We make this dedication for the benefit of the public at
-- large and to the detriment of our heirs and successors. We intend this 
-- dedication to be an overt act of relinquishment in perpetuity of all present
-- and future rights to this software under copyright law.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR 
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, 
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN 
-- ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION
-- WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
--
-- THIS DISCLAIMER MUST BE RETAINED AS PART OF THIS FILE AT ALL TIMES. 
-------------------------------------------------------------------------------

library work;
use work.esistream_pkg.all;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library STD;
use STD.textio.all;

library unisim;
use unisim.vcomponents.all;

entity tb_rx_esistream_top is
end entity tb_rx_esistream_top;

architecture behavioral of tb_rx_esistream_top is
---------------- Constants ----------------
  constant GEN_ESISTREAM       : boolean                               := true;
  constant GEN_GPIO            : boolean                               := true;
  constant NB_LANES            : natural                               := 8;
  constant COMMA               : std_logic_vector(31 downto 0)         := x"FF0000FF";
  signal sso_p                 : std_logic                             := '0';
  signal sso_n                 : std_logic                             := '1';
  signal FABRIC_CLK_P          : std_logic                             := '0';
  signal FABRIC_CLK_N          : std_logic                             := '1';
  signal clk_100mhz            : std_logic                             := '0';
  signal fmc_xcvr_out_p        : std_logic_vector(NB_LANES-1 downto 0) := (others => '0');
  signal fmc_xcvr_out_n        : std_logic_vector(NB_LANES-1 downto 0) := (others => '1');
  signal SW_C                  : std_logic                             := '0';
  signal SW_S                  : std_logic                             := '0';
  signal SW_W                  : std_logic                             := '0';
  signal SW_E                  : std_logic                             := '0';
  signal SW_N                  : std_logic                             := '0';
  signal dipswitch             : std_logic                             := '0';
  signal led_usr               : std_logic_vector(7 downto 0)          := (others => '0');
  --
  signal led_uart_ready        : std_logic                             := '0';
  signal led_sync_in           : std_logic                             := '0';
  signal led_ip_ready          : std_logic                             := '0';
  signal led_lanes_ready       : std_logic                             := '0';
  signal led_isrunning         : std_logic                             := '0';
  signal led_ber_status        : std_logic                             := '0';
  signal led_cb_status         : std_logic                             := '0';
  --
  signal tx_ip_ready           : std_logic                             := '0';
  signal rx_ip_ready           : std_logic                             := '0';
  signal ip_ready              : std_logic                             := '0';
  signal rx_lanes_ready        : std_logic                             := '0';
  signal tx_d_ctrl             : std_logic_vector(1 downto 0)          := (others => '0');
  signal pll_external_en       : std_logic                             := '0';
  signal rx_prbs_en            : std_logic                             := '0';
  signal tx_prbs_en            : std_logic                             := '0';
  signal tx_disp_en            : std_logic                             := '0';
  signal tx_lss                : std_logic                             := '0';
  signal start_stop_event      : std_logic                             := '0';
  signal change_data_mode      : std_logic                             := '0';
  signal sync                  : std_logic                             := '0';
  signal rst                   : std_logic                             := '0';
  signal rstn                  : std_logic                             := '0';
  signal rst_check             : std_logic                             := '0';
  signal ber_status            : std_logic                             := '0';
  signal cb_status             : std_logic                             := '0';
  constant STATUS_SUCCESS      : std_logic                             := '1';
  --
  signal aq600_rstn            : std_logic                             := '0';
  signal aq600_spi_sclk        : std_logic                             := '0';
  signal aq600_spi_csn         : std_logic                             := '0';
  signal LMX2592_CSN           : std_logic                             := '0';
  signal aq600_spi_mosi        : std_logic                             := '0';
  signal aq600_spi_miso        : std_logic                             := '0';
  signal PLL_LOCK              : std_logic                             := '0';
  signal aq600_synco_p         : std_logic                             := '0';
  signal aq600_synco_n         : std_logic                             := '0';
  signal aq600_synctrig_p      : std_logic                             := '0';
  signal aq600_synctrig_n      : std_logic                             := '0';
  --
  signal ASLp                  : std_logic_vector(1 downto 0)          := (others => '0');
  signal ASLn                  : std_logic_vector(1 downto 0)          := (others => '0');
  signal BSLp                  : std_logic_vector(1 downto 0)          := (others => '0');
  signal BSLn                  : std_logic_vector(1 downto 0)          := (others => '0');
  signal CSLp                  : std_logic_vector(1 downto 0)          := (others => '0');
  signal CSLn                  : std_logic_vector(1 downto 0)          := (others => '0');
  signal DSLp                  : std_logic_vector(1 downto 0)          := (others => '0');
  signal DSLn                  : std_logic_vector(1 downto 0)          := (others => '0');
--
  signal lfsr_init             : slv_17_array_n(NB_LANES-1 downto 0)   := (others => (others => '1'));
  signal clk_bit               : std_logic                             := '0';
  signal tx_clk                : std_logic                             := '0';
  signal txp                   : std_logic_vector(NB_LANES-1 downto 0) := (others => '0');
  signal txn                   : std_logic_vector(NB_LANES-1 downto 0) := (others => '1');
  constant NB_CLK_CYC          : std_logic_vector(31 downto 0)         := (others => '0');
  constant RST_CNTR_INIT       : std_logic_vector(11 downto 0)         := (others => '0');
  signal uart_tx               : std_logic                             := '0';
  signal uart_rx               : std_logic                             := '0';
  --
  -- -- UART IP constants:
  constant ADDR_RX_FIFO        : std_logic_vector(3 downto 0)          := x"0";
  constant ADDR_TX_FIFO        : std_logic_vector(3 downto 0)          := x"4";
  constant ADDR_STAT           : std_logic_vector(3 downto 0)          := x"8";
  constant ADDR_CTRL           : std_logic_vector(3 downto 0)          := x"C";
  --
  signal m1_axi_addr           : std_logic_vector(3 downto 0)          := (others => '0');
  signal m1_axi_strb           : std_logic_vector(3 downto 0)          := (others => '0');
  signal m1_axi_wdata          : std_logic_vector(31 downto 0)         := (others => '0');
  signal m1_axi_rdata          : std_logic_vector(31 downto 0)         := (others => '0');
  signal m1_axi_wen            : std_logic                             := '0';
  signal m1_axi_ren            : std_logic                             := '0';
  signal m1_axi_busy           : std_logic                             := '0';
  signal s1_interrupt          : std_logic                             := '0';
--
  signal reg_0_0, reg_0_1      : std_logic                             := '0';
  --
  signal reg3                  : std_logic_vector(7 downto 0)          := (others => '0');
  constant SPI_START_ENABLE    : std_logic_vector(7 downto 0)          := x"02";
  constant SPI_START_DISABLE   : std_logic_vector(7 downto 0)          := x"FD";
  constant SPI_SS_EXTERNAL_PLL : std_logic_vector(7 downto 0)          := x"01";
  constant SPI_SS_EV12AQ600    : std_logic_vector(7 downto 0)          := x"00";

begin
--
--############################################################################################################################
--############################################################################################################################
-- Clock Generation
--############################################################################################################################
--############################################################################################################################
  --sso_p  <= not sso_p  after 2.5 ns;
  --sso_n  <= not sso_n  after 2.5 ns;
  --
  FABRIC_CLK_P <= not FABRIC_CLK_P after 2.5 ns;
  FABRIC_CLK_N <= not FABRIC_CLK_N after 2.5 ns;
  --
  clk_100mhz   <= not clk_100mhz   after 5 ns;
  --
--############################################################################################################################
--############################################################################################################################
-- Unit under test
--############################################################################################################################
--############################################################################################################################   
  rx_esistream_top_1 : entity work.rx_esistream_top
    generic map (
      GEN_ESISTREAM          => GEN_ESISTREAM,
      GEN_GPIO               => GEN_GPIO,
      NB_LANES               => NB_LANES,
      RST_CNTR_INIT          => RST_CNTR_INIT,
      NB_CLK_CYC             => NB_CLK_CYC,
      CLK_MHz                => 100.0,
      SPI_CLK_MHz            => 10.0,
      SYNCTRIG_PULSE_WIDTH   => 7,
      SYNCTRIG_MAX_DELAY     => 10,
      SYNCTRIG_COUNTER_WIDTH => 8)
    port map (
      sso_n            => sso_n,
      sso_p            => sso_p,
      FABRIC_CLK_P     => FABRIC_CLK_P,
      FABRIC_CLK_N     => FABRIC_CLK_N,
      rxp              => txp,
      rxn              => txn,
      --ASLp             => ASLp,
      --ASLn             => ASLn,
      --BSLp             => BSLp,
      --BSLn             => BSLn,
      --CSLp             => CSLp,
      --CSLn             => CSLn,
      --DSLp             => DSLp,
      --DSLn             => DSLn,
      gpio_j20_10      => SW_C,
      gpio_j20_8       => SW_S,
      gpio_j20_6       => SW_W,
      gpio_j20_4       => SW_N,
      gpio_j20_2       => dipswitch,
      led_usr          => led_usr,
      UART_TX          => uart_tx,
      UART_RX          => uart_rx,
      aq600_rstn       => aq600_rstn,
      spi_sclk         => aq600_spi_sclk,
      spi_csn          => aq600_spi_csn,
      CSN_PLL          => LMX2592_CSN,
      spi_mosi         => aq600_spi_mosi,
      spi_miso         => aq600_spi_miso,
      PLL_LOCK         => PLL_LOCK,
      aq600_synco_p    => aq600_synco_p,
      aq600_synco_n    => aq600_synco_n,
      aq600_synctrig_p => aq600_synctrig_p,
      aq600_synctrig_n => aq600_synctrig_n);

  --ASLp(0)         <= txp(0);
  --ASLn(0)         <= txn(0);
  --ASLp(1)         <= txp(1);
  --ASLn(1)         <= txn(1);
  --BSLp(0)         <= txp(2);
  --BSLn(0)         <= txn(2);
  --BSLp(1)         <= txp(3);
  --BSLn(1)         <= txn(3);
  --CSLp(0)         <= txp(4);
  --CSLn(0)         <= txn(4);
  --CSLp(1)         <= txp(5);
  --CSLn(1)         <= txn(5);
  --DSLp(0)         <= txp(6);
  --DSLn(0)         <= txn(6);
  --DSLp(1)         <= txp(7);
  --DSLn(1)         <= txn(7);
  -- --
  dipswitch       <= rx_prbs_en;
  SW_C            <= rst;
  SW_S            <= sync;
  SW_W            <= rst_check;
  SW_N            <= '0';
  -- --
  led_uart_ready  <= led_usr(0);
  led_ip_ready    <= led_usr(1);
  led_lanes_ready <= led_usr(2);
  led_ber_status  <= led_usr(3);
  led_cb_status   <= led_usr(4);
  -- <= led_usr(6);
  reg_0_0         <= led_usr(6);
  reg_0_1         <= led_usr(7);
  --
  rx_ip_ready     <= led_ip_ready;
  ip_ready        <= tx_ip_ready and rx_ip_ready;
--============================================================================================================================
-- Stimulus
--============================================================================================================================
  my_tb : process
    -- 
    procedure axi4_lite_write
      (
        signal clk         : in  std_logic;
        constant addr      : in  std_logic_vector;
        constant data      : in  std_logic_vector;
        signal m_axi_addr  : out std_logic_vector;
        signal m_axi_strb  : out std_logic_vector;
        signal m_axi_wdata : out std_logic_vector;
        signal m_axi_wen   : out std_logic;
        signal m_axi_busy  : in  std_logic) is
    begin
      wait until rising_edge(clk);
      m_axi_addr  <= addr;
      m_axi_strb  <= "0001";
      m_axi_wdata <= x"000000"&data;
      m_axi_wen   <= '1';
      wait until rising_edge(clk);
      m_axi_wen   <= '0';
      wait until falling_edge(m_axi_busy);
    end axi4_lite_write;
    --
    procedure axi4_lite_read
      (
        signal clk         : in  std_logic;
        constant addr      : in  std_logic_vector;
        signal rdata       : out std_logic_vector;
        signal m_axi_addr  : out std_logic_vector;
        signal m_axi_rdata : in  std_logic_vector;
        signal m_axi_ren   : out std_logic;
        signal m_axi_busy  : in  std_logic) is
    begin
      wait until rising_edge(clk);
      m_axi_addr <= addr;
      m_axi_ren  <= '1';
      wait until rising_edge(clk);
      m_axi_ren  <= '0';
      wait until falling_edge(m_axi_busy);
      rdata      <= m_axi_rdata;
    end axi4_lite_read;
  begin
    -------------------------------- 
    -- tb init
    -------------------------------- 
    rst        <= '1';
    rst_check  <= '1';
    rx_prbs_en <= '1';
    tx_prbs_en <= '1';
    tx_disp_en <= '1';
    tx_d_ctrl  <= "01";  -- [01 : positive ramp mode]
    reg3       <= SPI_SS_EV12AQ600;
    --reg3     <= SPI_SS_EXTERNAL_PLL;
    sync       <= '0';
    wait for 100 ns;
    rst_check  <= '0';
    wait for 100 ns;
    rst        <= '0';
    report "start testbench... release reset.";
    ----------------------------------------------------------------------------------------------------
    -- TEST 1: 
    ---------------------------------------------------------------------------------------------------- 
    wait for 1000 ns;
    wait until rising_edge(clk_100mhz);
    rst        <= '1';
    wait until rising_edge(clk_100mhz);
    rst        <= '0';

    wait until rising_edge(led_ip_ready);
    wait for 100 ns;
    wait until rising_edge(clk_100mhz);
    sync <= '1';
    wait until rising_edge(clk_100mhz);
    sync <= '0';

    wait until rising_edge(led_lanes_ready);    
    wait for 100 ns;
    rst_check  <= '1';
    wait for 100 ns;
    rst_check  <= '0';
    ----------------------------------------------------------------------------------------------------
    -- TEST 2: Comment TEST 1 and set boolean constant GEN_ESISTREAM to false to speed up simulation for
    -- uart & spi communication tests below.
    -- uart 115200, 8-bit
    ----------------------------------------------------------------------------------------------------
    report "start testbench... release reset.";
    wait until rising_edge(led_uart_ready);
    -------------------------------- 
    -- s1 enable interrupt of tb uart_wrapper_1 module
    -------------------------------- 
    axi4_lite_write(clk_100mhz, ADDR_CTRL, x"10", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);  -- s1 enable interrupt
    wait for 200 us;

    -------------------------------- 
    -- UART WRITE command 
    --------------------------------
    -- spi slave select command, external pll
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"00", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"03", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"00", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"00", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"00", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, reg3, m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    wait for 1 ms;
    wait until rising_edge(clk_100mhz);
    -- spi write fifo in 
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"00", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"04", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"00", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"55", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"AA", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"55", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    wait for 1 ms;
    wait until rising_edge(clk_100mhz);
    -- spi write fifo in 
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"00", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"04", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"00", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"87", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"65", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"43", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    --
    reg3 <= reg3 or SPI_START_ENABLE;
    wait for 1 ms;
    wait until rising_edge(clk_100mhz);
    -- spi start command
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"00", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"03", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"00", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"00", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, x"00", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    axi4_lite_write(clk_100mhz, ADDR_TX_FIFO, reg3, m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);
    wait for 1 ms;
    wait until rising_edge(clk_100mhz);
    -- wait until rising_edge(s1_interrupt);                                                                     -- Wait TX FIFO empty
    -- wait until rising_edge(s1_interrupt);                                                                     -- Wait ACK
    -- axi4_lite_read(clk, ADDR_RX_FIFO, s1_rdata, m1_axi_addr, m1_axi_rdata, m1_axi_ren, m1_axi_busy);
    -- -- axi4_lite_write(clk_100mhz, ADDR_CTRL, x"10", m1_axi_addr, m1_axi_strb, m1_axi_wdata, m1_axi_wen, m1_axi_busy);  -- s1 enable interrupt
    -- -- wait until rising_edge(s1_interrupt);                                                                     -- Wait TX FIFO empty
    -- -- wait until rising_edge(s1_interrupt);                                                                     -- Wait ACK
    -- -- axi4_lite_read(clk_100mhz, ADDR_RX_FIFO, s1_rdata, m1_axi_addr, m1_axi_rdata, m1_axi_ren, m1_axi_busy);
    assert false report "Test finish" severity failure;
    wait;
  end process;

  gen_esistream_hdl : if GEN_ESISTREAM = true generate
    -- esistream clock generation:
    --clk_bit <= not clk_bit after 40.0 ps;    -- KU060 min clk bit period 80 ps
    --clk_bit <= not clk_bit after 39.0625 ps; -- KU040 
    clk_bit <= not clk_bit after 50.0 ps;      -- 7VX690

    tx_esistream_emulator_1 : entity work.tx_emu_esistream_top
      generic map (
        NB_LANES => NB_LANES,
        COMMA    => COMMA)
      port map (
        rst         => rst,
        clk         => clk_bit,
        sync_in     => aq600_synctrig_p,
        prbs_en     => tx_prbs_en,
        disp_en     => tx_disp_en,
        lfsr_init   => lfsr_init,
        data_ctrl   => tx_d_ctrl,
        sso_p       => sso_p,
        sso_n       => sso_n,
        tx_clk      => tx_clk,
        tx_ip_ready => tx_ip_ready,
        txp         => txp,
        txn         => txn,
        lss         => tx_lss);  -- when '1' lane synchronization sequence (FAS + PSS) sent on txp/n lanes else normal data.
  end generate gen_esistream_hdl;

  -- Simulate PC:
  rstn <= not rst;
  uart_wrapper_1 : entity work.uart_wrapper
    port map (
      clk         => clk_100mhz,
      rstn        => rstn,
      m_axi_addr  => m1_axi_addr,
      m_axi_strb  => m1_axi_strb,
      m_axi_wdata => m1_axi_wdata,
      m_axi_rdata => m1_axi_rdata,
      m_axi_wen   => m1_axi_wen,
      m_axi_ren   => m1_axi_ren,
      m_axi_busy  => m1_axi_busy,
      interrupt   => s1_interrupt,
      tx          => uart_tx,
      rx          => uart_rx);
--
end behavioral;
